library verilog;
use verilog.vl_types.all;
entity tbench is
end tbench;
